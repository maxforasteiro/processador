module instruction_data(clock, instruction_address, instruction_data_output);
  input clock;
  input [31:0] instruction_address;
  output [31:0] instruction_data_output;
  reg [31:0] instruction_ram [40:0];
  integer first_load = 0;
  
  always @ (posedge clock) begin
    if(first_load == 0) begin
		instruction_ram[0] = 32'b00100_000000000000000000000000000;
		instruction_ram[1] = 32'b01011_11101_00000_00000000000000001;
		instruction_ram[2] = 32'b01100_11110_0000000000000000000000;
		instruction_ram[3] = 32'b01101_11110_0000000000000000000000;
		instruction_ram[4] = 32'b00100_000000000000000000000000000;
		instruction_ram[5] = 32'b00111_11110_11101_00000000000011001;
		
		//##PROG 1##
		instruction_ram[6] = 32'b01011_00001_00000_00000000000000000;
		instruction_ram[7] = 32'b01011_00010_00000_00000000000000001;
		instruction_ram[8] = 32'b01100_00011_0000000000000000000000;
		instruction_ram[9] = 32'b01101_00011_0000000000000000000000;
		instruction_ram[10] = 32'b00100_000000000000000000000000000;
		instruction_ram[11] = 32'b01011_00100_00000_00000000000000001;
		instruction_ram[12] = 32'b01011_01010_00000_00000000000000000;
		instruction_ram[13] = 32'b00000_00010_00001_01010000000000000;
		instruction_ram[14] = 32'b00001_00001_00010_00000000000000000;
		instruction_ram[15] = 32'b00001_00010_01010_00000000000000000;
		instruction_ram[16] = 32'b00001_00100_00100_00000000000000001;
		instruction_ram[17] = 32'b01101_00010_0000000000000000000000;
		instruction_ram[18] = 32'b00100_000000000000000000000000000;
		instruction_ram[19] = 32'b01000_00100_00011_00000000000001101;
		instruction_ram[20] = 32'b00100_000000000000000000000000000;
		instruction_ram[21] = 32'b01101_00010_0000000000000000000000;
		instruction_ram[22] = 32'b01110_00010_00000_00000000000000001;
		instruction_ram[23] = 32'b00101_000000000000000000000000000;
		instruction_ram[24] = 32'b00110_00000_0000000000000000000000;
		
		
		//##PROG 2
		instruction_ram[25] = 32'b01011_00001_00000_00000000000000011;
		instruction_ram[26] = 32'b01011_00010_00000_00000000000000111;
		instruction_ram[27] = 32'b01111_00001_00010_00011000000000000;
		instruction_ram[28] = 32'b00010_00010_00011_00100000000000000;
		instruction_ram[29] = 32'b01101_00100_0000000000000000000000;
		instruction_ram[30] = 32'b01010_01010_00000_00000000000000001;
		instruction_ram[31] = 32'b01001_01010_00000_00101_000000000000;
		instruction_ram[32] = 32'b01101_00101_0000000000000000000000;
		instruction_ram[33] = 32'b01011_00110_00000_00000000000001000;
		instruction_ram[34] = 32'b10001_00001_00110_01011000000000000;
		instruction_ram[35] = 32'b01101_01011_0000000000000000000000;
		instruction_ram[36] = 32'b01100_10100_0000000000000000000000;
		instruction_ram[37] = 32'b10110_00000_10100_10110_00010_00000_00;
		instruction_ram[38] = 32'b01101_10110_0000000000000000000000;
		instruction_ram[39] = 32'b00101_000000000000000000000000000;
		instruction_ram[40] = 32'b00110_00000_0000000000000000000000;
		first_load = 1;
    end
  end
  
  assign instruction_data_output = instruction_ram[instruction_address];
endmodule