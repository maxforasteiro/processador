library verilog;
use verilog.vl_types.all;
entity extende_to_reg_size_vlg_vec_tst is
end extende_to_reg_size_vlg_vec_tst;
