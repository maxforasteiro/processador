library verilog;
use verilog.vl_types.all;
entity processing_unit_vlg_vec_tst is
end processing_unit_vlg_vec_tst;
