library verilog;
use verilog.vl_types.all;
entity mux_4_vlg_vec_tst is
end mux_4_vlg_vec_tst;
