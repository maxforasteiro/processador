library verilog;
use verilog.vl_types.all;
entity register_base_vlg_vec_tst is
end register_base_vlg_vec_tst;
