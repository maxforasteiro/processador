library verilog;
use verilog.vl_types.all;
entity instruction_data_vlg_vec_tst is
end instruction_data_vlg_vec_tst;
