library verilog;
use verilog.vl_types.all;
entity program_counter_vlg_vec_tst is
end program_counter_vlg_vec_tst;
