library verilog;
use verilog.vl_types.all;
entity ALUmodule_vlg_vec_tst is
end ALUmodule_vlg_vec_tst;
