library verilog;
use verilog.vl_types.all;
entity memory_data_vlg_vec_tst is
end memory_data_vlg_vec_tst;
