library verilog;
use verilog.vl_types.all;
entity ALU_module_vlg_vec_tst is
end ALU_module_vlg_vec_tst;
