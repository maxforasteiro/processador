library verilog;
use verilog.vl_types.all;
entity extender_vlg_vec_tst is
end extender_vlg_vec_tst;
