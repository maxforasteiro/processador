library verilog;
use verilog.vl_types.all;
entity extender_vlg_check_tst is
    port(
        extended        : in     vl_logic_vector(31 downto 0);
        sampler_rx      : in     vl_logic
    );
end extender_vlg_check_tst;
